module gateway

// Current API/Gateway Version
// fixme: move to a better location
pub const API_VERSION = "9"
