module gateway

// todo move out of gateway

pub enum OP_CODES {
	Dispatch
	Heartbeat
	Identify
	Presence_Update
	Voice_State_Update
	Resume
	Reconnect
	Request_Guild_Members
	Invalid_Session
	Hello
	Heartbeat_ACK
}

pub enum CLOSE_EVENT_CODES {
	UNKNOWN_ERROR = 4000
	UNKNOWN_OPCODE
	DECODE_ERROR
	NOT_AUTHENTICATED
	AUTHENTICATION_FAILED
	ALREADY_AUTHENTICATED
	INVALID_SEQ
	RATE_LIMITED
	SESSION_TIMED_OUT
	INVALID_SHARD
	SHARDING_REQUIRED
	INVALID_API_VERSION
	INVALID_INTENTS
	DISALLOWED_INTENTS
}

[flag]
pub enum GATEWAY_INTENTS {
	GUILDS = 1

	GUILD_MEMBERS = 1 << 1

	GUILD_BANS = 1 << 2

	GUILD_EMOJIS_AND_STICKERS = 1 << 3

	GUILD_INTEGRATIONS = 1 << 4

	GUILD_WEBHOOKS = 1 << 5

	GUILD_INVITES = 1 << 6

	GUILD_VOICE_STATES = 1 << 7

	GUILD_PRESENCES = 1 << 8

	GUILD_MESSAGES = 1 << 9

	GUILD_MESSAGE_REACTIONS = 1 << 10

	GUILD_MESSAGE_TYPING = 1 << 11

	DIRECT_MESSAGES = 1 << 12

	DIRECT_MESSAGE_REACTIONS = 1 << 13

	GUILD_SCHEDULED_EVENTS = 1 << 16
}
