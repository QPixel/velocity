module http


